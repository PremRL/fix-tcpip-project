----------------------------------------------------------------------------------
----------------------------------------------------------------------------------
-- Filename     Rom1024x8.vhd
-- Title        ROM for preparing FIX messages 
-- 
-- Author       L.Ratchanon
-- Date         2021/02/12
-- Syntax       VHDL
-- Remark       New Creation
-- Description    
--
----------------------------------------------------------------------------------
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
USE STD.TEXTIO.ALL;

Entity Rom1024x8 Is
	Port 
	(
		Clk			: in	std_logic;

		RdAddr		: in 	std_logic_vector( 9 downto 0);
		RdData		: out 	std_logic_vector( 7 downto 0)
	);
End Entity Rom1024x8;

Architecture rtl Of Rom1024x8 Is

----------------------------------------------------------------------------------
-- Constant declaration
----------------------------------------------------------------------------------
	
	constant ROM_DEPTH : integer := 1024;
	constant ROM_WIDTH : integer := 8;

	type array1024ofu8 is array (0 to ROM_DEPTH - 1) of std_logic_vector( ROM_WIDTH-1 downto 0);
	
	-- Notation 
	-- Each Market data content has 12 bytes
	-- First byte: 4 MSB is the address' distance for indexing frist symbol data 
	-- and 4 LSB is the address' distance for indexing frist SecurityID data 
	-- Next 6 byte: Storing Symbol of the corresponding market data 
	-- Last 5 byte: Storing SecurityID of the corresponding market data 	
	Constant ROMDATA 			: array1024ofu8 := 
		( x"12", x"41", x"44", x"56", x"41", x"4e", x"43", x"30", x"31", x"30", x"36", x"39", 
		  x"42", x"30", x"30", x"30", x"41", x"4f", x"54", x"30", x"31", x"31", x"31", x"37", 
		  x"41", x"30", x"30", x"30", x"41", x"57", x"43", x"34", x"36", x"38", x"34", x"36", 
		  x"42", x"30", x"30", x"30", x"42", x"42", x"4c", x"00", x"31", x"32", x"31", x"33", 
		  x"32", x"30", x"30", x"42", x"44", x"4d", x"53", x"00", x"31", x"32", x"31", x"39", 
		  x"41", x"30", x"30", x"30", x"42", x"45", x"4d", x"31", x"37", x"37", x"30", x"35", 
		  x"21", x"30", x"42", x"47", x"52", x"49", x"4d", x"32", x"37", x"34", x"30", x"33", 
		  x"52", x"30", x"30", x"30", x"30", x"42", x"48", x"30", x"31", x"32", x"32", x"32", 
		  x"42", x"30", x"30", x"30", x"42", x"4a", x"43", x"30", x"31", x"32", x"32", x"38", 
		  x"41", x"30", x"30", x"30", x"42", x"50", x"50", x"32", x"32", x"33", x"35", x"36", 
		  x"42", x"30", x"30", x"30", x"42", x"54", x"53", x"30", x"32", x"36", x"38", x"35", 
		  x"41", x"30", x"30", x"30", x"43", x"42", x"47", x"31", x"31", x"34", x"39", x"30", 
		  x"22", x"30", x"43", x"50", x"41", x"4c", x"4c", x"30", x"31", x"38", x"36", x"30", 
		  x"42", x"30", x"30", x"30", x"43", x"50", x"46", x"30", x"31", x"34", x"37", x"35", 
		  x"42", x"30", x"30", x"30", x"43", x"50", x"4e", x"30", x"31", x"34", x"39", x"39", 
		  x"41", x"30", x"30", x"30", x"43", x"52", x"43", x"35", x"31", x"30", x"33", x"36", 
		  x"32", x"30", x"30", x"44", x"54", x"41", x"43", x"30", x"31", x"38", x"33", x"31", 
		  x"52", x"30", x"30", x"30", x"30", x"45", x"41", x"30", x"35", x"34", x"34", x"35", 
		  x"32", x"30", x"30", x"45", x"47", x"43", x"4f", x"30", x"31", x"37", x"36", x"37", 
		  x"12", x"47", x"4c", x"4f", x"42", x"41", x"4c", x"30", x"32", x"36", x"33", x"38", 
		  x"31", x"30", x"30", x"47", x"50", x"53", x"43", x"31", x"33", x"39", x"37", x"39", 
		  x"31", x"30", x"30", x"47", x"55", x"4c", x"46", x"33", x"30", x"30", x"33", x"37", 
		  x"22", x"30", x"48", x"4d", x"50", x"52", x"4f", x"30", x"31", x"36", x"34", x"35", 
		  x"12", x"49", x"4e", x"54", x"55", x"43", x"48", x"30", x"32", x"37", x"39", x"35", 
		  x"32", x"30", x"30", x"49", x"52", x"50", x"43", x"30", x"31", x"37", x"31", x"31", 
		  x"42", x"30", x"30", x"30", x"49", x"56", x"4c", x"30", x"32", x"36", x"37", x"38", 
		  x"22", x"30", x"4b", x"42", x"41", x"4e", x"4b", x"30", x"31", x"38", x"31", x"37", 
		  x"42", x"30", x"30", x"30", x"4b", x"54", x"42", x"30", x"31", x"37", x"39", x"33", 
		  x"42", x"30", x"30", x"30", x"4b", x"54", x"43", x"30", x"31", x"38", x"31", x"34", 
		  x"52", x"30", x"30", x"30", x"30", x"4c", x"48", x"30", x"31", x"39", x"30", x"33", 
		  x"32", x"30", x"30", x"4d", x"49", x"4e", x"54", x"30", x"31", x"32", x"37", x"37", 
		  x"41", x"30", x"30", x"30", x"4d", x"54", x"43", x"31", x"31", x"35", x"38", x"38", 
		  x"41", x"30", x"30", x"30", x"4f", x"53", x"50", x"33", x"37", x"32", x"34", x"39", 
		  x"42", x"30", x"30", x"30", x"50", x"54", x"54", x"30", x"32", x"30", x"39", x"39", 
		  x"22", x"30", x"50", x"54", x"54", x"45", x"50", x"30", x"32", x"30", x"38", x"31", 
		  x"22", x"30", x"50", x"54", x"54", x"47", x"43", x"30", x"32", x"38", x"39", x"30", 
		  x"22", x"30", x"52", x"41", x"54", x"43", x"48", x"30", x"32", x"31", x"34", x"39", 
		  x"22", x"30", x"53", x"41", x"57", x"41", x"44", x"30", x"38", x"38", x"37", x"39", 
		  x"42", x"30", x"30", x"30", x"53", x"43", x"42", x"30", x"32", x"31", x"37", x"30", 
		  x"42", x"30", x"30", x"30", x"53", x"43", x"43", x"30", x"32", x"31", x"37", x"33", 
		  x"32", x"30", x"30", x"54", x"43", x"41", x"50", x"30", x"31", x"36", x"32", x"32", 
		  x"22", x"30", x"54", x"49", x"53", x"43", x"4f", x"30", x"32", x"35", x"36", x"32", 
		  x"42", x"30", x"30", x"30", x"54", x"4d", x"42", x"30", x"32", x"33", x"36", x"36", 
		  x"41", x"30", x"30", x"30", x"54", x"4f", x"41", x"32", x"39", x"32", x"32", x"30", 
		  x"42", x"30", x"30", x"30", x"54", x"4f", x"50", x"30", x"31", x"31", x"35", x"30", 
		  x"32", x"30", x"30", x"54", x"52", x"55", x"45", x"30", x"32", x"34", x"39", x"33", 
		  x"42", x"30", x"30", x"30", x"54", x"54", x"57", x"30", x"31", x"33", x"38", x"37", 
		  x"42", x"30", x"30", x"30", x"54", x"56", x"4f", x"30", x"32", x"34", x"32", x"32", 
		  x"42", x"30", x"30", x"30", x"56", x"47", x"49", x"30", x"34", x"39", x"35", x"39", 
		  x"21", x"30", x"57", x"48", x"41", x"55", x"50", x"32", x"35", x"35", x"36", x"33", 
		  -- 49 ROW Passing 
		  -- NOT USED 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  -- 59
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  -- 69
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  -- 79
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
		  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		  x"00", x"00", x"00", x"00" );
		  
----------------------------------------------------------------------------------
-- Signal declaration
----------------------------------------------------------------------------------
	
	signal rRdData				: std_logic_vector( 7 downto 0 );

Begin 
----------------------------------------------------------------------------------
-- Output assignment
----------------------------------------------------------------------------------
	
	RdData	<= rRdData;		
	
----------------------------------------------------------------------------------
-- DFF 
----------------------------------------------------------------------------------
	
	u_rRdData : Process (Clk) Is 
	Begin 
		if ( rising_edge(Clk) ) then 
			rRdData	<= ROMDATA(conv_integer(RdAddr));
		end if;
	End Process u_rRdData;

End Architecture rtl;